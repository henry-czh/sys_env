module core(
  input clk,
  input rst_n
);

initial begin
	$display("This is core Model!");
end

endmodule
